`ifndef WAVES
`define WAVES 8
`define SELECT_WIDTH $clog2(`WAVES)
`define WAVE_WIDTH 8
`define RANGE 32.0
`define range 32
`define max ((2**(`WAVE_WIDTH))-1)
`define MAX 255.0
`endif
