`ifndef WAVES
`define WAVES 8
`define SELECT_WIDTH $clog2(`WAVES)
`define WAVE_WIDTH 8
`endif
